library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 9
	
	
    );
   port (
          Endereco : in std_logic_vector (8 DOWNTO 0);
          Dado : out std_logic_vector (15 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0)   := "0000";
  constant LDA  : std_logic_vector(3 downto 0)   := "0001";
  constant SOMA : std_logic_vector(3 downto 0)   := "0010";
  constant SUB  : std_logic_vector(3 downto 0)   := "0011";
  constant LDI  : std_logic_vector(3 downto 0)   := "0100";
  constant STA  : std_logic_vector(3 downto 0)   := "0101";
  constant JMP	 : std_logic_vector(3 downto 0)   := "0110";
  constant JEQ  : std_logic_vector(3 downto 0)   := "0111";
  constant CEQ  : std_logic_vector(3 downto 0)   := "1000";
  constant JSR  : std_logic_vector(3 downto 0)   := "1001";
  constant RET  : std_logic_vector(3 downto 0)   := "1010";
  constant ANDOP  : std_logic_vector(3 downto 0) := "1011";
  constant CLT 	: std_logic_vector(3 downto 0) := "1100";
  constant JLT  : std_logic_vector(3 downto 0)   := "1101";
  
  -- Registradores
  
  constant RUS : std_logic_vector(2 downto 0) := "000"; -- Valor da unidade de segundos
  constant RDS : std_logic_vector(2 downto 0) := "001"; -- Valor da dezena de segundos
  constant RUM : std_logic_vector(2 downto 0) := "010"; -- Valor da unidade de minutos
  constant RDM : std_logic_vector(2 downto 0) := "011"; -- Valor da dezena de minutos
  constant RUH : std_logic_vector(2 downto 0) := "100"; -- Valor da unidade de horas
  constant RDH : std_logic_vector(2 downto 0) := "101"; -- Valor da dezena de horas
  
  constant RCA : std_logic_vector(2 downto 0) := "110"; -- Registrador para operaçoes aritméticas
  constant RCZ : std_logic_vector(2 downto 0) := "111"; -- Registrador de comparação com zero 


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  
-- INICIALIZACAO

--tmp(0)  := RCA & JSR & "000000010";  
--tmp(1)  := JMP & "000101001";  
--tmp(2)  := STA & "111111111";      -- Reseta o KEY0 
--tmp(3)  := STA & "111111110";      -- Reseta o KEY 1 
--tmp(4)  := LDI & "000000000";  
--tmp(5)  := STA & "000000000";      -- Constante 0 
--tmp(6)  := LDI & "000000001";  
--tmp(7)  := STA & "000000001";      -- Constante 1 
--tmp(8)  := LDI & "000001010";  
--tmp(9)  := STA & "000001010";      -- Constante 10 
--tmp(10)  := LDI & "000001001";  
--tmp(11)  := STA & "000001001";      -- Constante 9 
--tmp(12)  := LDI & "000001111";      -- Constante 15 : Mascara para SW 
--tmp(13)  := STA & "000001011";  
--tmp(14)  := LDA & "000000000";      -- Carrega o acumulador com o valor 0 
--tmp(15)  := STA & "100100000";      -- Limpa HEX0 
--tmp(16)  := STA & "100100001";      -- Limpa HEX1 
--tmp(17)  := STA & "100100010";      -- Limpa HEX2 
--tmp(18)  := STA & "100100011";      -- Limpa HEX3 
--tmp(19)  := STA & "100100100";      -- Limpa HEX4 
--tmp(20)  := STA & "100100101";      -- Limpa HEX5 
--tmp(21)  := STA & "100000000";      -- Limpa LEDR0~LEDR7 
--tmp(22)  := STA & "100000001";      -- Limpa LEDR8 
--tmp(23)  := STA & "100000010";      -- Limpa LEDR9 
--tmp(24)  := STA & "000000010";      -- Inicializa o Valor das unidades 
--tmp(25)  := STA & "000000011";      -- Inicializa o Valor das dezenas 
--tmp(26)  := STA & "000000100";      -- Inicializa o Valor das centenas 
--tmp(27)  := STA & "000000101";      -- Inicializa o Valor das unidade de milhares 
--tmp(28)  := STA & "000000110";      -- Inicializa o Valor das dezenas de milhares 
--tmp(29)  := STA & "000000111";      -- Inicializa o Valor das centenas de milhares 
--tmp(30)  := LDI & "000001010";  
--tmp(31)  := STA & "000001101";      -- Limite para o Valor das unidades 
--tmp(32)  := STA & "000001110";      -- Limite para o Valor das dezenas 
--tmp(33)  := STA & "000001111";      -- Limite para o Valor das centenas 
--tmp(34)  := STA & "000010000";      -- Limite para o Valor das unidade de milhares 
--tmp(35)  := STA & "000010001";      -- Limite para o Valor das dezenas de milhares 
--tmp(36)  := STA & "000010010";      -- Limite para o Valor das centenas de milhares 
--tmp(37)  := LDI & "000000000";  
--tmp(38)  := STA & "000001000";      -- Limpa a Flag de limite 
--tmp(39)  := STA & "000001100";      -- Limpa a Flag de Overflow(carry_out) 
--tmp(40)  := RET & "000000000";
--
--
--
---- LOOP_INICIO
--
--
--tmp(41)  := LDA & "101100000";      -- Carrega o acumulador com a leitura do botão KEY0 
--tmp(42)  := ANDOP & "000000001";  
--tmp(43)  := CEQ & "000000001";      -- Compara a leitura de KEY0 com a constante 1 MEM[1] 
--tmp(44)  := JEQ & "000111000";  
--tmp(45)  := JSR & "001111110";  
--tmp(46)  := LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
--tmp(47)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(48)  := CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
--tmp(49)  := JEQ & "000111100";  
--tmp(50)  := JSR & "010010111";  
--tmp(51)  := LDA & "101100100";      -- Carrega o acumulador com a leitura do botão FPGA_RESET 
--tmp(52)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(53)  := CEQ & "000000001";      -- Compara a leitura de FPGA_RESET com a constante 1 MEM[1] 
--tmp(54)  := JEQ & "000111010";  
--tmp(55)  := JMP & "000101001";  
--
--
---- INCREMENTA_CONTADOR_CHECKPOINT:
--
--
--tmp(56)  := JSR & "000111110";  
--tmp(57)  := JMP & "000101101";
--
--
---- REINICIA_CONTADOR_CHECKPOINT:
--
--
--tmp(58)  := JSR & "010001011";  
--tmp(59)  := JMP & "000110111"; 
--
---- LIMITE_INCREMENTO_CHECKPOINT:
--
--
--tmp(60)  := JSR & "010101101";  
--tmp(61)  := JMP & "000110010";
--
--
---- INCREMENTA_CONTADOR
--
--
--tmp(62)  := STA & "111111111";  
--tmp(63)  := LDA & "000001100";  
--tmp(64)  := CEQ & "000000001";  
--tmp(65)  := JEQ & "001111101";      -- Verifica o carry_out 
--tmp(66)  := LDA & "000001000";  
--tmp(67)  := CEQ & "000000001";  
--tmp(68)  := JEQ & "001111101";      -- Verifica o carry_out 
--tmp(69)  := LDA & "000000010";  
--tmp(70)  := SOMA & "000000001";  
--tmp(71)  := CEQ & "000001010";  
--tmp(72)  := JEQ & "001001011";      -- Verifica as unidades 
--tmp(73)  := STA & "000000010";  
--tmp(74)  := JMP & "001111101";  
--tmp(75)  := LDI & "000000000";  
--tmp(76)  := STA & "000000010";  
--tmp(77)  := LDA & "000000011";  
--tmp(78)  := SOMA & "000000001";  
--tmp(79)  := CEQ & "000001010";  
--tmp(80)  := JEQ & "001010011";      -- Verifica as dezenas 
--tmp(81)  := STA & "000000011";  
--tmp(82)  := JMP & "001111101";  
--tmp(83)  := LDI & "000000000";  
--tmp(84)  := STA & "000000011";  
--tmp(85)  := LDA & "000000100";  
--tmp(86)  := SOMA & "000000001";  
--tmp(87)  := CEQ & "000001010";  
--tmp(88)  := JEQ & "001011011";      -- Verifica as centenas 
--tmp(89)  := STA & "000000100";  
--tmp(90)  := JMP & "001111101";  
--tmp(91)  := LDI & "000000000";  
--tmp(92)  := STA & "000000100";  
--tmp(93)  := LDA & "000000101";  
--tmp(94)  := SOMA & "000000001";  
--tmp(95)  := CEQ & "000001010";  
--tmp(96)  := JEQ & "001100011";      -- Verifica as Unidade de Milhares 
--tmp(97)  := STA & "000000101";  
--tmp(98)  := JMP & "001111101";  
--tmp(99)  := LDI & "000000000";  
--tmp(100)  := STA & "000000101";  
--tmp(101)  := LDA & "000000110";  
--tmp(102)  := SOMA & "000000001";  
--tmp(103)  := CEQ & "000001010";  
--tmp(104)  := JEQ & "001101011";      -- Verifica as dezenas de Milhares 
--tmp(105)  := STA & "000000110";  
--tmp(106)  := JMP & "001111101";  
--tmp(107)  := LDI & "000000000";  
--tmp(108)  := STA & "000000110";  
--tmp(109)  := LDA & "000000111";  
--tmp(110)  := SOMA & "000000001";  
--tmp(111)  := CEQ & "000001010";  
--tmp(112)  := JEQ & "001110011";      -- Verifica as centenas de Milhares 
--tmp(113)  := STA & "000000111";  
--tmp(114)  := JMP & "001111101";  
--tmp(115)  := LDI & "000000001";  
--tmp(116)  := STA & "100000010";      -- Ativa o LED de OVERLFOW 
--tmp(117)  := STA & "000001100";      -- Ativa a Flag de OVERFLOW 
--tmp(118)  := LDI & "000001001";  
--tmp(119)  := STA & "000000010";      -- Mantem os valore das unidades em 9 
--tmp(120)  := STA & "000000011";      -- Mantem os valore das dezenas em 9 
--tmp(121)  := STA & "000000100";      -- Mantem os valore das centenas em 9 
--tmp(122)  := STA & "000000101";      -- Mantem os valore das unidades de milhares em 9 
--tmp(123)  := STA & "000000110";      -- Mantem os valore das dezenas de milhares em 9 
--tmp(124)  := STA & "000000111";      -- Mantem os valore das centenas de milhares em 9 
--tmp(125)  := RET & "000000000";  
--
---- ESCREVE_DISPLAY
--
--
--tmp(126)  := LDA & "000000010";  
--tmp(127)  := STA & "100100000";      -- Escreve o valor das unidades 
--tmp(128)  := LDA & "000000011";  
--tmp(129)  := STA & "100100001";      -- Escreve o valor das dezenas 
--tmp(130)  := LDA & "000000100";  
--tmp(131)  := STA & "100100010";      -- Escreve o valor das centenas 
--tmp(132)  := LDA & "000000101";  
--tmp(133)  := STA & "100100011";      -- Escreve o valor das unidades de milhares 
--tmp(134)  := LDA & "000000110";  
--tmp(135)  := STA & "100100100";      -- Escreve o valor das dezenas de milhares 
--tmp(136)  := LDA & "000000111";  
--tmp(137)  := STA & "100100101";      -- Escreve o valor das centenas de milhares 
--tmp(138)  := RET & "000000000";  
--
---- REINICIA_CONTADOR
--
--
--tmp(139)  := LDI & "000000000";  
--tmp(140)  := STA & "000000010";      -- Reinicia o Valor das unidades 
--tmp(141)  := STA & "000000011";      -- Reinicia o Valor das dezenas 
--tmp(142)  := STA & "000000100";      -- Reinicia o Valor das centenas 
--tmp(143)  := STA & "000000101";      -- Reinicia o Valor das unidade de milhares 
--tmp(144)  := STA & "000000110";      -- Reinicia o Valor das dezenas de milhares 
--tmp(145)  := STA & "000000111";      -- Reinicia o Valor das centenas de milhares 
--tmp(146)  := STA & "000001000";      -- Reinicia a Flag de Limite 
--tmp(147)  := STA & "000001100";      -- Reinicia a Falg de Overflow(carry_out) 
--tmp(148)  := STA & "100000001";      -- Apaga o Led de Limite 
--tmp(149)  := STA & "100000010";      -- Apaga o Led de Overflow 
--tmp(150)  := RET & "000000000"; 
--
--
---- VERIFICA_LIMITE
--
--
--tmp(151)  := LDA & "000000010";  
--tmp(152)  := CLT & "000001101";  
--tmp(153)  := JLT & "010101100";      -- Verifica as unidades 
--tmp(154)  := LDA & "000000011";  
--tmp(155)  := CLT & "000001110";  
--tmp(156)  := JLT & "010101100";      -- Verifica as dezenas 
--tmp(157)  := LDA & "000000100";  
--tmp(158)  := CLT & "000001111";  
--tmp(159)  := JLT & "010101100";      -- Verifica as centenas 
--tmp(160)  := LDA & "000000101";  
--tmp(161)  := CLT & "000010000";  
--tmp(162)  := JLT & "010101100";      -- Verifica as unidades de milhares 
--tmp(163)  := LDA & "000000110";  
--tmp(164)  := CLT & "000010001";  
--tmp(165)  := JLT & "010101100";      -- Verifica as dezenas de milhares 
--tmp(166)  := LDA & "000000111";  
--tmp(167)  := CLT & "000010010";  
--tmp(168)  := JLT & "010101100";      -- Verifica as centenas de milhares 
--tmp(169)  := LDI & "000000001";  
--tmp(170)  := STA & "000001000";      -- Flag de Limite 
--tmp(171)  := STA & "100000001";      -- LED de Limite 
--tmp(172)  := RET & "000000000";
--
--
---- LIMITE_INCREMENTO
--
--
--tmp(173)  := STA & "111111110";      -- Limpa a leitura do KEY1 
--tmp(174)  := LDI & "000000001";  
--tmp(175)  := STA & "100000000";      -- Liga o LEDR0 
--tmp(176)  := LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
--tmp(177)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(178)  := CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
--tmp(179)  := JEQ & "010111100";  
--tmp(180)  := LDA & "101000000";      -- Leitura SW 
--tmp(181)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(182)  := CLT & "000001010";  
--tmp(183)  := JLT & "010111010";  
--tmp(184)  := LDI & "000001001";  
--tmp(185)  := STA & "100100000";  
--tmp(186)  := STA & "100100000";  
--tmp(187)  := JMP & "010110000";  
--tmp(188)  := LDA & "101000000";      -- Leitura SW 
--tmp(189)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(190)  := CLT & "000001010";  
--tmp(191)  := JLT & "011000010";  
--tmp(192)  := LDI & "000001001";  
--tmp(193)  := STA & "000001101";      -- Guarda o Limite das unidades 
--tmp(194)  := STA & "000001101";  
--tmp(195)  := STA & "111111110";      -- Limpa a leitura do KEY1 
--tmp(196)  := LDI & "000000010";  
--tmp(197)  := STA & "100000000";      -- Liga o LEDR1 
--tmp(198)  := LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
--tmp(199)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(200)  := CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
--tmp(201)  := JEQ & "011010010";  
--tmp(202)  := LDA & "101000000";      -- Leitura SW 
--tmp(203)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(204)  := CLT & "000001010";  
--tmp(205)  := JLT & "011010000";  
--tmp(206)  := LDI & "000001001";  
--tmp(207)  := STA & "100100001";  
--tmp(208)  := STA & "100100001";  
--tmp(209)  := JMP & "011000110";  
--tmp(210)  := LDA & "101000000";      -- Leitura SW 
--tmp(211)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(212)  := CLT & "000001010";  
--tmp(213)  := JLT & "011011000";  
--tmp(214)  := LDI & "000001001";  
--tmp(215)  := STA & "000001110";      -- Guarda o Limite das dezenas 
--tmp(216)  := STA & "000001110";  
--tmp(217)  := STA & "111111110";      -- Limpa a leitura do KEY1 
--tmp(218)  := LDI & "000000100";  
--tmp(219)  := STA & "100000000";      -- Liga o LEDR2 
--tmp(220)  := LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
--tmp(221)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(222)  := CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
--tmp(223)  := JEQ & "011101000";  
--tmp(224)  := LDA & "101000000";      -- Leitura SW 
--tmp(225)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(226)  := CLT & "000001010";  
--tmp(227)  := JLT & "011100110";  
--tmp(228)  := LDI & "000001001";  
--tmp(229)  := STA & "100100010";  
--tmp(230)  := STA & "100100010";  
--tmp(231)  := JMP & "011011100";  
--tmp(232)  := LDA & "101000000";      -- Leitura SW 
--tmp(233)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(234)  := CLT & "000001010";  
--tmp(235)  := JLT & "011101110";  
--tmp(236)  := LDI & "000001001";  
--tmp(237)  := STA & "000001111";      -- Guarda o Limite das centenas 
--tmp(238)  := STA & "000001111";  
--tmp(239)  := STA & "111111110";      -- Limpa a leitura do KEY1 
--tmp(240)  := LDI & "000001000";  
--tmp(241)  := STA & "100000000";      -- Liga o LEDR3 
--tmp(242)  := LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
--tmp(243)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(244)  := CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
--tmp(245)  := JEQ & "011111110";  
--tmp(246)  := LDA & "101000000";      -- Leitura SW 
--tmp(247)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(248)  := CLT & "000001010";  
--tmp(249)  := JLT & "011111100";  
--tmp(250)  := LDI & "000001001";  
--tmp(251)  := STA & "100100011";  
--tmp(252)  := STA & "100100011";  
--tmp(253)  := JMP & "011110010";  
--tmp(254)  := LDA & "101000000";      -- Leitura SW 
--tmp(255)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(256)  := CLT & "000001010";  
--tmp(257)  := JLT & "100000100";  
--tmp(258)  := LDI & "000001001";  
--tmp(259)  := STA & "000010000";      -- Guarda o Limite das unidade de milhares 
--tmp(260)  := STA & "000010000";  
--tmp(261)  := STA & "111111110";      -- Limpa a leitura do KEY1 
--tmp(262)  := LDI & "000010000";  
--tmp(263)  := STA & "100000000";      -- Liga o LEDR4 
--tmp(264)  := LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
--tmp(265)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(266)  := CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
--tmp(267)  := JEQ & "100010100";  
--tmp(268)  := LDA & "101000000";      -- Leitura SW 
--tmp(269)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(270)  := CLT & "000001010";  
--tmp(271)  := JLT & "100010010";  
--tmp(272)  := LDI & "000001001";  
--tmp(273)  := STA & "100100100";  
--tmp(274)  := STA & "100100100";  
--tmp(275)  := JMP & "100001000";  
--tmp(276)  := LDA & "101000000";      -- Leitura SW 
--tmp(277)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(278)  := CLT & "000001010";  
--tmp(279)  := JLT & "100011010";  
--tmp(280)  := LDI & "000001001";  
--tmp(281)  := STA & "000010001";      -- Guarda o Limite das dezenas de milhares 
--tmp(282)  := STA & "000010001";  
--tmp(283)  := STA & "111111110";      -- Limpa a leitura do KEY1 
--tmp(284)  := LDI & "000100000";  
--tmp(285)  := STA & "100000000";      -- Liga o LEDR5 
--tmp(286)  := LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
--tmp(287)  := ANDOP & "000000001";      -- Aplica mascara 
--tmp(288)  := CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
--tmp(289)  := JEQ & "100101010";  
--tmp(290)  := LDA & "101000000";      -- Leitura SW 
--tmp(291)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(292)  := CLT & "000001010";  
--tmp(293)  := JLT & "100101000";  
--tmp(294)  := LDI & "000001001";  
--tmp(295)  := STA & "100100101";  
--tmp(296)  := STA & "100100101";  
--tmp(297)  := JMP & "100011110";  
--tmp(298)  := LDA & "101000000";      -- Leitura SW 
--tmp(299)  := ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
--tmp(300)  := CLT & "000001010";  
--tmp(301)  := JLT & "100110000";  
--tmp(302)  := LDI & "000001001";  
--tmp(303)  := STA & "000010010";      -- Guarda o Limite das centenas de milhares 
--tmp(304)  := STA & "000010010";  
--tmp(305)  := LDI & "000000000";  
--tmp(306)  := STA & "100100000";      -- Limpa o HEX0 
--tmp(307)  := STA & "100100001";      -- Limpa o HEX1 
--tmp(308)  := STA & "100100001";      -- Limpa o HEX2 
--tmp(309)  := STA & "100100010";      -- Limpa o HEX3 
--tmp(310)  := STA & "100100011";      -- Limpa o HEX4 
--tmp(311)  := STA & "100000000";      -- Limpa o HEX5 
--tmp(312)  := STA & "111111110";      -- Limpa a leitura do KEY1 
--tmp(313)  := RET & "000000000";  
--return tmp;
tmp(0)  := RCA & JSR & "000000010";  
tmp(1)  := RCA & JMP & "000110001";  
tmp(2)  := RCZ & LDI & "000000000";      -- Registrador com zero 
tmp(3)  := RCZ & STA & "111111111";      -- Reseta o KEY0 
tmp(4)  := RCZ & STA & "111111110";      -- Reseta o KEY 1 
tmp(5)  := RCZ & STA & "000000000";      -- Constante 0 
tmp(6)  := RCA & LDI & "000000001";  
tmp(7)  := RCA & STA & "000000001";      -- Constante 1 
tmp(8)  := RCA & LDI & "000000010";      -- Constante 2 
tmp(9)  := RCA & STA & "000000010";  
tmp(10)  := RCA & LDI & "000000011";      -- Constante 3 
tmp(11)  := RCA & STA & "000000011";  
tmp(12)  := RCA & LDI & "000000100";      -- Constante 4 
tmp(13)  := RCA & STA & "000000100";  
tmp(14)  := RCA & LDI & "000000110";      -- Constante 6 
tmp(15)  := RCA & STA & "000000110";  
tmp(16)  := RCA & LDI & "000001010";  
tmp(17)  := RCA & STA & "000001010";      -- Constante 10 
tmp(18)  := RCA & LDI & "000001001";  
tmp(19)  := RCA & STA & "000001001";      -- Constante 9 
tmp(20)  := RCA & LDI & "000001111";      -- Constante 15 : Mascara para SW 
tmp(21)  := RCA & STA & "000001011";  
tmp(22)  := RCZ & STA & "100100000";      -- Limpa HEX0 
tmp(23)  := RCZ & STA & "100100001";      -- Limpa HEX1 
tmp(24)  := RCZ & STA & "100100010";      -- Limpa HEX2 
tmp(25)  := RCZ & STA & "100100011";      -- Limpa HEX3 
tmp(26)  := RCZ & STA & "100100100";      -- Limpa HEX4 
tmp(27)  := RCZ & STA & "100100101";      -- Limpa HEX5 
tmp(28)  := RCZ & STA & "100000000";      -- Limpa LEDR0~LEDR7 
tmp(29)  := RCZ & STA & "100000001";      -- Limpa LEDR8 
tmp(30)  := RCZ & STA & "100000010";      -- Limpa LEDR9 
tmp(31)  := RUS & LDI & "000000000";      -- Inicializa o Valor das unidades de segundos 
tmp(32)  := RDS & LDI & "000000000";      -- Inicializa o Valor das dezenas de segundos 
tmp(33)  := RUM & LDI & "000000000";      -- Inicializa o Valor das unidades de minutos 
tmp(34)  := RDM & LDI & "000000000";      -- Inicializa o Valor das dezenas de minutos 
tmp(35)  := RUH & LDI & "000000000";      -- Inicializa o Valor das unidades de horas 
tmp(36)  := RDH & LDI & "000000000";      -- Inicializa o Valor das dezenas de horas 
tmp(37)  := RCA & LDI & "000001010";  
tmp(38)  := RCA & STA & "000001101";      -- Limite para o Valor das unidades de segundos 
tmp(39)  := RCA & STA & "000001110";      -- Limite para o Valor das dezenas de segundos 
tmp(40)  := RCA & STA & "000001111";      -- Limite para o Valor das unidades de minutos 
tmp(41)  := RCA & STA & "000010000";      -- Limite para o Valor das dezenas de minutos 
tmp(42)  := RCA & STA & "000010001";      -- Limite para o Valor das unidades de horas 
tmp(43)  := RCA & STA & "000010010";      -- Limite para o Valor das dezenas de horas 
tmp(44)  := RCZ & STA & "000001000";      -- Limpa a Flag de limite 
tmp(45)  := RCZ & STA & "000001100";      -- Limpa a Flag de Overflow(carry_out) 
tmp(46)  := RCZ & STA & "000011011";      -- Inicializa o valor para lidar com formato de hora 
tmp(47)  := RCZ & STA & "000011100";      -- Inicializa o valor para lidar com limite de 24 Horas 
tmp(48)  := RCZ & RET & "000000000";  
tmp(49)  := RCA & LDA & "101100000";      -- Carrega o acumulador com a leitura do botão KEY0 
tmp(50)  := RCA & ANDOP & "000000001";  
tmp(51)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY0 com a constante 1 MEM[1] 
tmp(52)  := RCA & JEQ & "001000100";  
tmp(53)  := RCA & JSR & "010000011";  
tmp(54)  := RCA & LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(55)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(56)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(57)  := RCA & JEQ & "001001000";  
tmp(58)  := RCA & JSR & "010010110";  
tmp(59)  := RCA & LDA & "101100100";      -- Carrega o acumulador com a leitura do botão FPGA_RESET 
tmp(60)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(61)  := RCA & CEQ & "000000001";      -- Compara a leitura de FPGA_RESET com a constante 1 MEM[1] 
tmp(62)  := RCA & JEQ & "001000110";  
tmp(63)  := RCA & LDA & "101100010";      -- Carrega o acumulador com a leitura do botão KEY2 
tmp(64)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(65)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY2 com a constante 1 MEM[1] 
tmp(66)  := RCA & JEQ & "001001010";  
tmp(67)  := RCA & JMP & "000110001";  
tmp(68)  := RCA & JSR & "001001100";  
tmp(69)  := RCA & JMP & "000110101";  
tmp(70)  := RCA & JSR & "010001010";  
tmp(71)  := RCA & JMP & "000111111";  
tmp(72)  := RCA & JSR & "010100110";  
tmp(73)  := RCA & JMP & "000111010";  
tmp(74)  := RCA & JSR & "101001111";  
tmp(75)  := RCA & JMP & "001000011";  
tmp(76)  := RCA & STA & "111111111";  
tmp(77)  := RCA & LDA & "000001100";  
tmp(78)  := RCA & CEQ & "000000001";  
tmp(79)  := RCA & JEQ & "010000010";      -- Verifica o carry_out 
tmp(80)  := RCA & LDA & "000001000";  
tmp(81)  := RCA & CEQ & "000000001";  
tmp(82)  := RCA & JEQ & "010000010";      -- Verifica o carry_out 
tmp(83)  := RUS & SOMA & "000000001";  
tmp(84)  := RUS & CEQ & "000001010";  
tmp(85)  := RCA & JEQ & "001010111";      -- Verifica as unidades de segundos 
tmp(86)  := RCA & JMP & "010000010";  
tmp(87)  := RUS & LDI & "000000000";  
tmp(88)  := RDS & SOMA & "000000001";  
tmp(89)  := RDS & CEQ & "000000110";  
tmp(90)  := RCA & JEQ & "001011100";      -- Verifica as dezenas de segundos 
tmp(91)  := RCA & JMP & "010000010";  
tmp(92)  := RDS & LDI & "000000000";  
tmp(93)  := RUM & SOMA & "000000001";  
tmp(94)  := RUM & CEQ & "000001010";  
tmp(95)  := RCA & JEQ & "001100001";      -- Verifica as unidades de minutos 
tmp(96)  := RCA & JMP & "010000010";  
tmp(97)  := RUM & LDI & "000000000";  
tmp(98)  := RDM & SOMA & "000000001";  
tmp(99)  := RDM & CEQ & "000000110";  
tmp(100)  := RCA & JEQ & "001100110";      -- Verifica as dezenas de minutos 
tmp(101)  := RCA & JMP & "010000010";  
tmp(102)  := RDM & LDI & "000000000";  
tmp(103)  := RUH & SOMA & "000000001";  
tmp(104)  := RUH & CEQ & "000000100";  
tmp(105)  := RCA & JEQ & "001101011";  
tmp(106)  := RCA & JMP & "001110000";  
tmp(107)  := RCA & LDA & "000011011";  
tmp(108)  := RCA & SOMA & "000000001";  
tmp(109)  := RCA & STA & "000011011";  
tmp(110)  := RCA & CEQ & "000000011";  
tmp(111)  := RCA & JEQ & "001111000";  
tmp(112)  := RUH & CEQ & "000001010";  
tmp(113)  := RCA & JEQ & "001110011";      -- Verifica as unidades de horas 
tmp(114)  := RCA & JMP & "010000010";  
tmp(115)  := RUH & LDI & "000000000";  
tmp(116)  := RDH & SOMA & "000000001";  
tmp(117)  := RDH & CEQ & "000000011";  
tmp(118)  := RCA & JEQ & "001111000";      -- Verifica  a dezena das horas 
tmp(119)  := RCA & JMP & "010000010";  
tmp(120)  := RCA & LDI & "000000001";  
tmp(121)  := RCA & STA & "100000010";      -- Ativa o LED de OVERLFOW 
tmp(122)  := RCA & STA & "000001100";      -- Ativa a Flag de OVERFLOW 
tmp(123)  := RUS & LDI & "000001001";      -- Mantem os valore das unidades de segundos em 9 
tmp(124)  := RDS & LDI & "000000101";      -- Mantem os valore das dezenas de segundos 5 
tmp(125)  := RUM & LDI & "000001001";      -- Mantem os valore das unidades de minutos em 9 
tmp(126)  := RDM & LDI & "000000101";      -- Mantem os valore das dezenas de minutos em 5 
tmp(127)  := RUH & LDI & "000000011";      -- Mantem os valore das unidades de horas em 3 
tmp(128)  := RDH & LDI & "000000010";      -- Mantem os valore das dezenas em 2 
tmp(129)  := RCZ & STA & "000011011";  
tmp(130)  := RCZ & RET & "000000000";  
tmp(131)  := RUS & STA & "100100000";      -- Escreve o valor das unidades de segundos 
tmp(132)  := RDS & STA & "100100001";      -- Escreve o valor das dezenas de segundos 
tmp(133)  := RUM & STA & "100100010";      -- Escreve o valor das unidades de minutos 
tmp(134)  := RDM & STA & "100100011";      -- Escreve o valor das dezenas de minutos 
tmp(135)  := RUH & STA & "100100100";      -- Escreve o valor das unidades de horas 
tmp(136)  := RDH & STA & "100100101";      -- Escreve o valor das dezenas de horas 
tmp(137)  := RDH & RET & "000000000";  
tmp(138)  := RUS & LDI & "000000000";      -- Reinicia os valores das unidades de segundos em 9 
tmp(139)  := RDS & LDI & "000000000";      -- Renicia os valores das dezenas de segundos 5 
tmp(140)  := RUM & LDI & "000000000";      -- Reinicia os valores das unidades de minutos em 9 
tmp(141)  := RDM & LDI & "000000000";      -- Reinicia os valores das dezenas de minutos em 5 
tmp(142)  := RUH & LDI & "000000000";      -- Reinicia os valores das unidades de horas em 3 
tmp(143)  := RDH & LDI & "000000000";      -- Reinicia os valores das dezenas de horas em 2 
tmp(144)  := RCZ & STA & "000001000";      -- Reinicia a Flag de Limite 
tmp(145)  := RCZ & STA & "000001100";      -- Reinicia a Falg de Overflow(carry_out) 
tmp(146)  := RCZ & STA & "100000001";      -- Apaga o Led de Limite 
tmp(147)  := RCZ & STA & "100000010";      -- Apaga o Led de Overflow 
tmp(148)  := RCZ & STA & "000011011";      -- Reinicia a contagem de formato 24 
tmp(149)  := RCZ & RET & "000000000";  
tmp(150)  := RUS & CLT & "000001101";  
tmp(151)  := RCA & JLT & "010100101";      -- Verifica as unidades de segundos 
tmp(152)  := RDS & CLT & "000001110";  
tmp(153)  := RCA & JLT & "010100101";      -- Verifica as dezenas de segundos 
tmp(154)  := RUM & CLT & "000001111";  
tmp(155)  := RCA & JLT & "010100101";      -- Verifica as unidades de minutos 
tmp(156)  := RDM & CLT & "000010000";  
tmp(157)  := RCA & JLT & "010100101";      -- Verifica as dezenas de minutos 
tmp(158)  := RUH & CLT & "000010001";  
tmp(159)  := RCA & JLT & "010100101";      -- Verifica as unidades de horas 
tmp(160)  := RDH & CLT & "000010010";  
tmp(161)  := RCA & JLT & "010100101";      -- Verifica as dezenas de hpras 
tmp(162)  := RCA & LDI & "000000001";  
tmp(163)  := RCA & STA & "000001000";      -- Flag de Limite 
tmp(164)  := RCA & STA & "100000001";      -- LED de Limite 
tmp(165)  := RCA & RET & "000000000";  
tmp(166)  := RCZ & STA & "100100000";      -- Limpa HEX0 
tmp(167)  := RCZ & STA & "100100001";      -- Limpa HEX1 
tmp(168)  := RCZ & STA & "100100010";      -- Limpa HEX2 
tmp(169)  := RCZ & STA & "100100011";      -- Limpa HEX3 
tmp(170)  := RCZ & STA & "100100100";      -- Limpa HEX4 
tmp(171)  := RCZ & STA & "100100101";      -- Limpa HEX5 
tmp(172)  := RCZ & STA & "111111110";      -- Limpa a leitura do KEY1 
tmp(173)  := RCA & LDI & "000100000";  
tmp(174)  := RCA & STA & "100000000";      -- Liga o LEDR5 
tmp(175)  := RCA & LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(176)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(177)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(178)  := RCA & JEQ & "010111100";  
tmp(179)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(180)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(181)  := RCA & CLT & "000000011";  
tmp(182)  := RCA & JLT & "010111010";  
tmp(183)  := RCA & LDI & "000000001";  
tmp(184)  := RCA & STA & "000011100";  
tmp(185)  := RCA & LDI & "000000010";  
tmp(186)  := RCA & STA & "100100101";  
tmp(187)  := RCA & JMP & "010101111";  
tmp(188)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(189)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(190)  := RCA & CLT & "000000011";  
tmp(191)  := RCA & JLT & "011000011";  
tmp(192)  := RCA & LDI & "000000001";  
tmp(193)  := RCA & STA & "000011100";  
tmp(194)  := RCA & LDI & "000000010";      -- Guarda o Limite das dezenas de horas 
tmp(195)  := RCA & STA & "000010010";  
tmp(196)  := RCZ & STA & "111111110";      -- Limpa a leitura do KEY1 
tmp(197)  := RCA & LDI & "000010000";  
tmp(198)  := RCA & STA & "100000000";      -- Liga o LEDR4 
tmp(199)  := RCA & LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(200)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(201)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(202)  := RCA & JEQ & "011011110";  
tmp(203)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(204)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(205)  := RCA & LDA & "000011100";  
tmp(206)  := RCA & CEQ & "000000001";  
tmp(207)  := RCA & JEQ & "011010111";  
tmp(208)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(209)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(210)  := RCA & CLT & "000001010";  
tmp(211)  := RCA & JLT & "011011100";  
tmp(212)  := RCA & LDI & "000001001";  
tmp(213)  := RCA & STA & "100100100";  
tmp(214)  := RCA & JMP & "011011100";  
tmp(215)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(216)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(217)  := RCA & CLT & "000000100";  
tmp(218)  := RCA & JLT & "011011100";  
tmp(219)  := RCA & LDI & "000000011";  
tmp(220)  := RCA & STA & "100100100";  
tmp(221)  := RCA & JMP & "011000111";  
tmp(222)  := RCA & LDA & "000011100";  
tmp(223)  := RCA & CEQ & "000000001";  
tmp(224)  := RCA & JEQ & "011101000";  
tmp(225)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(226)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(227)  := RCA & CLT & "000001010";  
tmp(228)  := RCA & JLT & "011101101";  
tmp(229)  := RCA & LDI & "000001001";  
tmp(230)  := RCA & STA & "000010001";      -- Guarda o Limite das unidades de horas 
tmp(231)  := RCA & JMP & "011101101";  
tmp(232)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(233)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(234)  := RCA & CLT & "000000100";  
tmp(235)  := RCA & JLT & "011011100";  
tmp(236)  := RCA & LDI & "000000011";  
tmp(237)  := RCA & STA & "000010001";  
tmp(238)  := RCZ & STA & "111111110";      -- Limpa a leitura do KEY1 
tmp(239)  := RCA & LDI & "000001000";  
tmp(240)  := RCA & STA & "100000000";      -- Liga o LEDR3 
tmp(241)  := RCA & LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(242)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(243)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(244)  := RCA & JEQ & "011111101";  
tmp(245)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(246)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(247)  := RCA & CLT & "000000110";  
tmp(248)  := RCA & JLT & "011111011";  
tmp(249)  := RCA & LDI & "000000101";  
tmp(250)  := RCA & STA & "100100011";  
tmp(251)  := RCA & STA & "100100011";  
tmp(252)  := RCA & JMP & "011110001";  
tmp(253)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(254)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(255)  := RCA & CLT & "000000110";  
tmp(256)  := RCA & JLT & "100000011";  
tmp(257)  := RCA & LDI & "000000101";  
tmp(258)  := RCA & STA & "000010000";      -- Guarda o Limite das dezenas de minutos 
tmp(259)  := RCA & STA & "000010000";  
tmp(260)  := RCZ & STA & "111111110";      -- Limpa a leitura do KEY1 
tmp(261)  := RCA & LDI & "000000100";  
tmp(262)  := RCA & STA & "100000000";      -- Liga o LEDR2 
tmp(263)  := RCA & LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(264)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(265)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(266)  := RCA & JEQ & "100010011";  
tmp(267)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(268)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(269)  := RCA & CLT & "000001010";  
tmp(270)  := RCA & JLT & "100010001";  
tmp(271)  := RCA & LDI & "000001001";  
tmp(272)  := RCA & STA & "100100010";  
tmp(273)  := RCA & STA & "100100010";  
tmp(274)  := RCA & JMP & "100000111";  
tmp(275)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(276)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(277)  := RCA & CLT & "000001010";  
tmp(278)  := RCA & JLT & "100011001";  
tmp(279)  := RCA & LDI & "000001001";  
tmp(280)  := RCA & STA & "000001111";      -- Guarda o Limite das unidades de minutos 
tmp(281)  := RCA & STA & "000001111";  
tmp(282)  := RCZ & STA & "111111110";      -- Limpa a leitura do KEY1 
tmp(283)  := RCA & LDI & "000000010";  
tmp(284)  := RCA & STA & "100000000";      -- Liga o LEDR1 
tmp(285)  := RCA & LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(286)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(287)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(288)  := RCA & JEQ & "100101001";  
tmp(289)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(290)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(291)  := RCA & CLT & "000000110";  
tmp(292)  := RCA & JLT & "100100111";  
tmp(293)  := RCA & LDI & "000000101";  
tmp(294)  := RCA & STA & "100100001";  
tmp(295)  := RCA & STA & "100100001";  
tmp(296)  := RCA & JMP & "100011101";  
tmp(297)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(298)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(299)  := RCA & CLT & "000000110";  
tmp(300)  := RCA & JLT & "100101111";  
tmp(301)  := RCA & LDI & "000000101";  
tmp(302)  := RCA & STA & "000001110";      -- Guarda o Limite das dezenas de segundos 
tmp(303)  := RCA & STA & "000001110";  
tmp(304)  := RCZ & STA & "111111110";      -- Limpa a leitura do KEY1 
tmp(305)  := RCA & LDI & "000000001";  
tmp(306)  := RCA & STA & "100000000";      -- Liga o LEDR0 
tmp(307)  := RCA & LDA & "101100001";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(308)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(309)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(310)  := RCA & JEQ & "100111111";  
tmp(311)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(312)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(313)  := RCA & CLT & "000001010";  
tmp(314)  := RCA & JLT & "100111101";  
tmp(315)  := RCA & LDI & "000001001";  
tmp(316)  := RCA & STA & "100100000";  
tmp(317)  := RCA & STA & "100100000";  
tmp(318)  := RCA & JMP & "100110011";  
tmp(319)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(320)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(321)  := RCA & CLT & "000001010";  
tmp(322)  := RCA & JLT & "101000101";  
tmp(323)  := RCA & LDI & "000001001";  
tmp(324)  := RCA & STA & "000001101";      -- Guarda o Limite das unidades de segundos 
tmp(325)  := RCA & STA & "000001101";  
tmp(326)  := RCZ & STA & "100100000";      -- Limpa o HEX0 
tmp(327)  := RCZ & STA & "100100001";      -- Limpa o HEX1 
tmp(328)  := RCZ & STA & "100100001";      -- Limpa o HEX2 
tmp(329)  := RCZ & STA & "100100010";      -- Limpa o HEX3 
tmp(330)  := RCZ & STA & "100100011";      -- Limpa o HEX4 
tmp(331)  := RCZ & STA & "100000000";      -- Limpa o HEX5 
tmp(332)  := RCZ & STA & "111111110";      -- Limpa a leitura do KEY1 
tmp(333)  := RCZ & STA & "000011100";  
tmp(334)  := RCZ & RET & "000000000";  
tmp(335)  := RCZ & STA & "100100000";      -- Limpa HEX0 
tmp(336)  := RCZ & STA & "100100001";      -- Limpa HEX1 
tmp(337)  := RCZ & STA & "100100010";      -- Limpa HEX2 
tmp(338)  := RCZ & STA & "100100011";      -- Limpa HEX3 
tmp(339)  := RCZ & STA & "100100100";      -- Limpa HEX4 
tmp(340)  := RCZ & STA & "100100101";      -- Limpa HEX5 
tmp(341)  := RCZ & STA & "111111101";      -- Limpa a leitura do KEY2 
tmp(342)  := RCA & LDI & "000100000";  
tmp(343)  := RCA & STA & "100000000";      -- Liga o LEDR5 
tmp(344)  := RCA & LDA & "101100010";      -- Carrega o acumulador com a leitura do botão KEY2 
tmp(345)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(346)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(347)  := RCA & JEQ & "101100101";  
tmp(348)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(349)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(350)  := RCA & CLT & "000000011";  
tmp(351)  := RCA & JLT & "101100011";  
tmp(352)  := RCA & LDI & "000000001";  
tmp(353)  := RCA & STA & "000011100";  
tmp(354)  := RCA & LDI & "000000010";  
tmp(355)  := RCA & STA & "100100101";  
tmp(356)  := RCA & JMP & "101011000";  
tmp(357)  := RDH & LDA & "101000000";      -- Leitura SW 
tmp(358)  := RDH & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(359)  := RDH & CLT & "000000011";  
tmp(360)  := RCA & JLT & "101101100";  
tmp(361)  := RDH & LDI & "000000001";  
tmp(362)  := RDH & STA & "000011100";  
tmp(363)  := RDH & LDI & "000000010";      -- Guarda o Limite das dezenas de horas 
tmp(364)  := RCZ & STA & "111111101";      -- Limpa a leitura do KEY2 
tmp(365)  := RCA & LDI & "000010000";  
tmp(366)  := RCA & STA & "100000000";      -- Liga o LEDR4 
tmp(367)  := RCA & LDA & "101100010";      -- Carrega o acumulador com a leitura do botão KEY1 
tmp(368)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(369)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(370)  := RCA & JEQ & "110000110";  
tmp(371)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(372)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(373)  := RCA & LDA & "000011100";  
tmp(374)  := RCA & CEQ & "000000001";  
tmp(375)  := RCA & JEQ & "101111111";  
tmp(376)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(377)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(378)  := RCA & CLT & "000001010";  
tmp(379)  := RCA & JLT & "110000100";  
tmp(380)  := RCA & LDI & "000001001";  
tmp(381)  := RCA & STA & "100100100";  
tmp(382)  := RCA & JMP & "110000100";  
tmp(383)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(384)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(385)  := RCA & CLT & "000000100";  
tmp(386)  := RCA & JLT & "110000100";  
tmp(387)  := RCA & LDI & "000000011";  
tmp(388)  := RCA & STA & "100100100";  
tmp(389)  := RCA & JMP & "101101111";  
tmp(390)  := RCA & LDA & "000011100";  
tmp(391)  := RCA & CEQ & "000000001";  
tmp(392)  := RCA & JEQ & "110001111";  
tmp(393)  := RUH & LDA & "101000000";      -- Leitura SW 
tmp(394)  := RUH & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(395)  := RUH & CLT & "000001010";  
tmp(396)  := RCA & JLT & "110010100";  
tmp(397)  := RUH & LDI & "000001001";  
tmp(398)  := RCA & JMP & "110010100";  
tmp(399)  := RUH & LDA & "101000000";      -- Leitura SW 
tmp(400)  := RUH & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(401)  := RUH & CLT & "000000100";  
tmp(402)  := RUH & JLT & "110000100";  
tmp(403)  := RUH & LDI & "000000011";  
tmp(404)  := RCZ & STA & "111111101";      -- Limpa a leitura do KEY2 
tmp(405)  := RCA & LDI & "000001000";  
tmp(406)  := RCA & STA & "100000000";      -- Liga o LEDR3 
tmp(407)  := RCA & LDA & "101100010";      -- Carrega o acumulador com a leitura do botão KEY2 
tmp(408)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(409)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(410)  := RCA & JEQ & "110100011";  
tmp(411)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(412)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(413)  := RCA & CLT & "000000110";  
tmp(414)  := RCA & JLT & "110100001";  
tmp(415)  := RCA & LDI & "000000101";  
tmp(416)  := RCA & STA & "100100011";  
tmp(417)  := RCA & STA & "100100011";  
tmp(418)  := RCA & JMP & "110010111";  
tmp(419)  := RDM & LDA & "101000000";      -- Leitura SW 
tmp(420)  := RDM & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(421)  := RDM & CLT & "000000110";  
tmp(422)  := RCA & JLT & "110101000";  
tmp(423)  := RDM & LDI & "000000101";  
tmp(424)  := RCZ & STA & "111111101";      -- Limpa a leitura do KEY2 
tmp(425)  := RCA & LDI & "000000100";  
tmp(426)  := RCA & STA & "100000000";      -- Liga o LEDR2 
tmp(427)  := RCA & LDA & "101100010";      -- Carrega o acumulador com a leitura do botão KEY2 
tmp(428)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(429)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(430)  := RCA & JEQ & "110110111";  
tmp(431)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(432)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(433)  := RCA & CLT & "000001010";  
tmp(434)  := RCA & JLT & "110110101";  
tmp(435)  := RCA & LDI & "000001001";  
tmp(436)  := RCA & STA & "100100010";  
tmp(437)  := RCA & STA & "100100010";  
tmp(438)  := RCA & JMP & "110101011";  
tmp(439)  := RUM & LDA & "101000000";      -- Leitura SW 
tmp(440)  := RUM & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(441)  := RUM & CLT & "000001010";  
tmp(442)  := RCA & JLT & "110111100";  
tmp(443)  := RUM & LDI & "000001001";  
tmp(444)  := RCZ & STA & "111111101";      -- Limpa a leitura do KEY2 
tmp(445)  := RCA & LDI & "000000010";  
tmp(446)  := RCA & STA & "100000000";      -- Liga o LEDR1 
tmp(447)  := RCA & LDA & "101100010";      -- Carrega o acumulador com a leitura do botão KEY2 
tmp(448)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(449)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(450)  := RCA & JEQ & "111001011";  
tmp(451)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(452)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(453)  := RCA & CLT & "000000110";  
tmp(454)  := RCA & JLT & "111001001";  
tmp(455)  := RCA & LDI & "000000101";  
tmp(456)  := RCA & STA & "100100001";  
tmp(457)  := RCA & STA & "100100001";  
tmp(458)  := RCA & JMP & "110111111";  
tmp(459)  := RDS & LDA & "101000000";      -- Leitura SW 
tmp(460)  := RDS & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(461)  := RDS & CLT & "000000110";  
tmp(462)  := RCA & JLT & "111010000";  
tmp(463)  := RDS & LDI & "000000101";  
tmp(464)  := RCZ & STA & "111111101";      -- Limpa a leitura do KEY2 
tmp(465)  := RCA & LDI & "000000001";  
tmp(466)  := RCA & STA & "100000000";      -- Liga o LEDR0 
tmp(467)  := RCA & LDA & "101100010";      -- Carrega o acumulador com a leitura do botão KEY2 
tmp(468)  := RCA & ANDOP & "000000001";      -- Aplica mascara 
tmp(469)  := RCA & CEQ & "000000001";      -- Compara a leitura de KEY1 com a constante 1 MEM[1] 
tmp(470)  := RCA & JEQ & "111011111";  
tmp(471)  := RCA & LDA & "101000000";      -- Leitura SW 
tmp(472)  := RCA & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(473)  := RCA & CLT & "000001010";  
tmp(474)  := RCA & JLT & "111011101";  
tmp(475)  := RCA & LDI & "000001001";  
tmp(476)  := RCA & STA & "100100000";  
tmp(477)  := RCA & STA & "100100000";  
tmp(478)  := RCA & JMP & "111010011";  
tmp(479)  := RUS & LDA & "101000000";      -- Leitura SW 
tmp(480)  := RUS & ANDOP & "000001011";      -- Aplica mascara SW0~SW3 
tmp(481)  := RUS & CLT & "000001010";  
tmp(482)  := RUS & JLT & "111100100";  
tmp(483)  := RUS & LDI & "000001001";  
tmp(484)  := RCZ & STA & "100100000";      -- Limpa o HEX0 
tmp(485)  := RCZ & STA & "100100001";      -- Limpa o HEX1 
tmp(486)  := RCZ & STA & "100100001";      -- Limpa o HEX2 
tmp(487)  := RCZ & STA & "100100010";      -- Limpa o HEX3 
tmp(488)  := RCZ & STA & "100100011";      -- Limpa o HEX4 
tmp(489)  := RCZ & STA & "100000000";      -- Limpa o HEX5 
tmp(490)  := RCZ & STA & "111111101";      -- Limpa a leitura do KEY1 
tmp(491)  := RCZ & STA & "000011100";  
tmp(492)  := RCZ & RET & "000000000";  
return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;